module divSig (output [19:0] m, input [9:0] a,b);
